-- This is the HyperRAM clock synthesis.
--
-- Created by Michael Jørgensen in 2022 (mjoergen.github.io/HyperRAM).

library ieee;
use ieee.std_logic_1164.all;

library unisim;
use unisim.vcomponents.all;

library xpm;
use xpm.vcomponents.all;

entity mega65_clk is
   port (
      sys_clk_i : in  std_logic;   -- expects 100 MHz
      sys_rst_i : in  std_logic;   -- Asynchronous, asserted low
      vga_clk_o : out std_logic;   -- 74.25 MHz
      vga_rst_o : out std_logic
   );
end entity mega65_clk;

architecture synthesis of mega65_clk is

   signal mmcm_fb   : std_logic;
   signal mmcm_clk  : std_logic;
   signal clk_fb    : std_logic;
   signal locked    : std_logic;

begin

   -- generate HyperRAM clock.
   -- VCO frequency range for Artix 7 speed grade -1 : 600 MHz - 1200 MHz
   -- f_VCO = f_CLKIN * CLKFBOUT_MULT_F / DIVCLK_DIVIDE   
   i_clk_mmcm : MMCME2_ADV
      generic map (
         BANDWIDTH            => "OPTIMIZED",
         CLKOUT4_CASCADE      => FALSE,
         COMPENSATION         => "ZHOLD",
         STARTUP_WAIT         => FALSE,
         CLKIN1_PERIOD        => 10.0,       -- INPUT @ 100 MHz
         REF_JITTER1          => 0.010,
         DIVCLK_DIVIDE        => 4,
         CLKFBOUT_MULT_F      => 37.125,
         CLKFBOUT_PHASE       => 0.000,
         CLKFBOUT_USE_FINE_PS => FALSE,
         CLKOUT0_DIVIDE_F     => 12.500,     -- 74.25 MHz
         CLKOUT0_PHASE        => 0.000,
         CLKOUT0_DUTY_CYCLE   => 0.500,
         CLKOUT0_USE_FINE_PS  => FALSE
      )
      port map (
         -- Output clocks
         CLKFBOUT            => mmcm_fb,
         CLKOUT0             => mmcm_clk,
         -- Input clock control
         CLKFBIN             => clk_fb,
         CLKIN1              => sys_clk_i,
         CLKIN2              => '0',
         -- Tied to always select the primary input clock
         CLKINSEL            => '1',
         -- Ports for dynamic reconfiguration
         DADDR               => (others => '0'),
         DCLK                => '0',
         DEN                 => '0',
         DI                  => (others => '0'),
         DO                  => open,
         DRDY                => open,
         DWE                 => '0',
         -- Ports for dynamic phase shift
         PSCLK               => '0',
         PSEN                => '0',
         PSINCDEC            => '0',
         PSDONE              => open,
         -- Other control and status signals
         LOCKED              => locked,
         CLKINSTOPPED        => open,
         CLKFBSTOPPED        => open,
         PWRDWN              => '0',
         RST                 => '0'
      ); -- i_clk_mmcm


   -------------------------------------
   -- Output buffering
   -------------------------------------

   i_bufg_clk_fb : BUFG
      port map (
         I => mmcm_fb,
         O => clk_fb
      ); -- i_bufg_clkfb

   i_bufg_clk : BUFG
      port map (
         I => mmcm_clk,
         O => vga_clk_o
      ); -- i_bufg_clk


   -------------------------------------
   -- Reset generation
   -------------------------------------

   i_xpm_cdc_sync_rst_pixel : xpm_cdc_sync_rst
      generic map (
         INIT_SYNC_FF => 1  -- Enable simulation init values
      )
      port map (
         src_rst  => not (not sys_rst_i and locked),  -- 1-bit input: Source reset signal.
         dest_clk => vga_clk_o,                       -- 1-bit input: Destination clock.
         dest_rst => vga_rst_o                        -- 1-bit output: src_rst synchronized to the destination clock domain.
                                                   -- This output is registered.
      ); -- i_xpm_cdc_sync_rst_pixel

end architecture synthesis;

